localparam RS =  552927 ;
