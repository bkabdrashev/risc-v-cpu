localparam RS =  507068 ;
